----------------------------------------------------------------------------------------------
-- Lab 5																												  --
-- ROM																												  --
-- Steve Comer																										  --
-- Edward Hazeldine																								  --
-- Michial Stikkel 																								  --
-- Updated 29 Oct 2012																							  --
-- 	Saves the Values in ROM																					  --
----------------------------------------------------------------------------------------------

-- Import the necessary libraries.
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

----------------------------------------------------------------------------------------------

ENTITY ROM IS

PORT(
	clk     : IN STD_LOGIC;
	address : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	dataOut : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);

END ROM;

ARCHITECTURE Behavioral OF ROM IS

	TYPE tROM IS ARRAY (0 TO 95) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
	CONSTANT cROM : tROM := (
--		-----------------------------------
--		-- TEST PROGRAM for CMPA, SUBA
--		0	=> "0000",  -- Load Acc
--		1  => "0101",	-- 	with 5
--		2  => "1001",	-- SUBAcc
--		3  => "0010",	--		with 2
--		4  => "1000",  -- ADDAcc
--		5  => "0011",	-- 	with 3
--		6	=> "1010",  -- CMPAcc
--		7  => "0110",	-- 	with 6, sets z flag
--		8  => "0011",	-- Display Acc
--		9  => "0110",	--		Displays 6
--		10 => "0000",	--
--		11 => "1010",  -- CMPAcc
--		12 => "1111",	-- 	with F
--		13 => "1000",  -- ADDAcc
--		14 => "0001",	-- 	with 1, turns off Z flag
--		15 => "0011",  -- Display Acc
--	   16 => "0110",	-- 	Displays 7
--		17 => "0000",  --
--		-----------------------------------
	
--		-----------------------------------
--		-- TEST PROGRAM for BEQ
--		0 	=> "0000",	-- Load Acc
--		1  => "0100",	--		with 4
--		2	=> "1000",	-- ADDAcc
--		3  => "0001",	-- 	with 1, Acc = 5
--		4	=> "1010",  -- CMPAcc
--		5  => "0101",	-- 	with 5
--		6  => "1100",	-- Branch if (Acc == 5)
--		7  => "0000",	--		to @0x02
--		8  => "0010",	--
--		9  => "0011",	-- Display Acc
--		10 => "0110",	--		Displays 6 if working
--		11 => "0000",	--		Displays 5 if BEQ doesn't work, 7 if BNE doesn't work
--		12 => "1010",	-- CMPAcc
--		13 => "0110",  -- 	with 6
--		14 => "1101",	-- Branch if (Acc != 6)
--		15 => "0000",	--		to @0x02
--		16 => "0010",	--
--		17	=> "1000",	-- ADDAcc
--		18 => "0001",	-- 	with 1
--		19 => "0011",	-- Display Acc
--		20 => "0110",	--		Displays 7 if working
--		21 => "0000",	--		Displays 8 if BEQ doesn't work
--		-----------------------------------

--		-----------------------------------
--		-- TEST PROGRAM for BEQ
--		0 	=> "0000",	-- loadA
--		1	=> "0011",	--    with 3
--		2	=> "0011",	-- store A
--		3	=> "1000",	-- @ 0x80
--		4  => "0000",	--
--		5 	=> "0000",	-- loadA
--		6	=> "0110",	--		with 6
--		7	=> "0011",	-- store A
--		8	=> "1000",	-- @ 0x81
--		9  => "0001",	--
--		10 => "0000",	-- loadA
--		11	=> "0000",	--		with 0
--		12	=> "0011",	-- store A
--		13	=> "1000",	-- @ 0x 82
--		14 => "0010",	--
--		15 => "0000",	-- loadA
--		16 => "0001",	-- 	with 1
--		17 => "1011",	-- BRA
--		18 => "1000",	-- to 0x80
--		19 => "0000",	--
--		-- Should display 1 to PORTLED from RAM
--		-- RAM 0x80 = 3
--		-- RAM 0x81 = 6
--		--	RAM 0x82 = 0
--		-- Displays 1 to PORTLED
--		-----------------------------------
		
		
		0  => "0000",
		1  => "0001",
		2  => "0011",
		3  => "0110",
		4  => "0000",
		5  => "1000",
		6  => "0010",
		7  => "0011",
		8  => "0110",
		9  => "0000",
		10 => "0110",
		11 => "0100",
		12 => "0101",
		13 => "1101",
		14 => "0011",
		15 => "0110",
		16 => "0000",
		17 => "1000",
		18 => "0011",
		19 => "0111",
		20 => "0011",
		21 => "0110",
		22 => "0000",
		23 => "1000",
		24 => "0010",
		25 => "1010",
		26 => "1111",
		27 => "1101",
		28 => "0001",
		29 => "0100",
		30 => "0011",
		31 => "0110",
------------------------------------	
		32 => "0000",
		33 => "1110",
		34 => "0010",
		35 => "0001",
		36 => "0100",
		37 => "0100",
		38 => "1000",
		39 => "0000",
		40 => "1111",
		41 => "1010",
		42 => "1110",
		43 => "1101",
		44 => "0010",
		45 => "0010",
		46 => "0001",
		47 => "0101",
		48 => "1110",
		49 => "0011",
		50 => "1000",
		51 => "0011",
		52 => "0001",
		53 => "0101",
		54 => "1111",
		55 => "0011",
		56 => "1000",
		57 => "0110",
		58 => "0000",
		59 => "1000",
		60 => "0011",
		61 => "1000",
		62 => "1000",
		63 => "1001",
------------------------------------
		64 => "1000",
		65 => "0011",
		66 => "1000",
		67 => "1001",
		68 => "0000",
		69 => "1011",
		70 => "0011",
		71 => "1000",
		72 => "1101",
		73 => "0000",
		74 => "0101",
		75 => "0011",
		76 => "1000",
		77 => "1110",
		78 => "0000",
		79 => "0110",
		80 => "0011",
		81 => "1000",
		82 => "1111",
		83 => "1011",
		84 => "1000",
		85 => "0000",
		86 => "1100",
		87 => "0000",
		88 => "0000",
		89 => "0000",
		90 => "1110",
		91 => "0011",
		92 => "0110",
		93 => "0000",
		94 => "1001",
		95 => "0000");
	 
BEGIN

	Read_Process : PROCESS(clk)	
	BEGIN
		IF rising_edge(clk) THEN
			dataOut <= cROM(conv_integer(address));
		END IF;
	END PROCESS Read_Process;
	
		
END Behavioral;